// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Sun Dec 22 20:02:10 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module location_sm (
    input wire reset,
    input wire clock,
    input wire station1,
    input wire station0,
    output reg [5:0] total_loc
	 );

    
    reg [10:0] fstate;
    reg [10:0] reg_fstate;
    parameter init=0,stable=1,st1=2,stable1=3,st2=4,stable2=5,st3=6,stable3=7,st4=8,stable4=9,st5=10;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or station1 or station0)
    begin
        if (reset) begin
            reg_fstate <= init;
            total_loc <= 6'b000000;
        end
        else begin
            total_loc <= 6'b000000;
            case (fstate)
                init: begin
                    if ((station1 == 1'b1))
                        reg_fstate <= stable;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= init;

                    total_loc <= 6'b000001;
                end
                stable: begin
                    if ((station0 == 1'b1))
                        reg_fstate <= st1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable;

                    total_loc <= 6'b000001;
                end
                st1: begin
                    if ((station0 == 1'b0))
                        reg_fstate <= stable1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st1;

                    total_loc <= 6'b000010;
                end
                stable1: begin
                    if ((station0 == 1'b1))
                        reg_fstate <= st2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable1;

                    total_loc <= 6'b000010;
                end
                st2: begin
                    if ((station0 == 1'b0))
                        reg_fstate <= stable2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st2;

                    total_loc <= 6'b000100;
                end
                stable2: begin
                    if ((station0 == 1'b1))
                        reg_fstate <= st3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable2;

                    total_loc <= 6'b000100;
                end
                st3: begin
                    if ((station0 == 1'b0))
                        reg_fstate <= stable3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st3;

                    total_loc <= 6'b001000;
                end
                stable3: begin
                    if ((station0 == 1'b1))
                        reg_fstate <= st4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable3;

                    total_loc <= 6'b001000;
                end
                st4: begin
                    if ((station0 == 1'b0))
                        reg_fstate <= stable4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st4;

                    total_loc <= 6'b010000;
                end
                stable4: begin
                    if ((station0 == 1'b1))
                        reg_fstate <= st5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable4;

                    total_loc <= 6'b010000;
                end
                st5: begin
                    if ((station0 == 1'b0))
                        reg_fstate <= st5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st5;

                    total_loc <= 6'b100000;
                end
                default: begin
                    total_loc <= 6'bxxxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // location_sm
