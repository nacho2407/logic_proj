// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Wed Dec 11 22:19:14 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module speed_control_sm (
    reset,clock,under_limit,cur_spd3,cur_spd2,cur_spd1,cur_spd0,tik,
    emerg_stop);

    input reset;
    input clock;
    input under_limit;
    input cur_spd3;
    input cur_spd2;
    input cur_spd1;
    input cur_spd0;
    input tik;
    tri0 reset;
    tri0 under_limit;
    tri0 cur_spd3;
    tri0 cur_spd2;
    tri0 cur_spd1;
    tri0 cur_spd0;
    tri0 tik;
    output emerg_stop;
    reg emerg_stop;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter stable=0,warning1=1,warning2=2,stop=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or under_limit or cur_spd3 or cur_spd2 or cur_spd1 or cur_spd0 or tik)
    begin
        if (reset) begin
            reg_fstate <= stable;
            emerg_stop <= 1'b0;
        end
        else begin
            emerg_stop <= 1'b0;
            case (fstate)
                stable: begin
                    if (((under_limit == 1'b0) & (tik == 1'b1)))
                        reg_fstate <= warning1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable;

                    emerg_stop <= 1'b0;
                end
                warning1: begin
                    if (((under_limit == 1'b0) & (tik == 1'b1)))
                        reg_fstate <= warning2;
                    else if ((under_limit == 1'b1))
                        reg_fstate <= stable;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= warning1;

                    emerg_stop <= 1'b0;
                end
                warning2: begin
                    if (((under_limit == 1'b0) & (tik == 1'b1)))
                        reg_fstate <= stop;
                    else if ((under_limit == 1'b1))
                        reg_fstate <= stable;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= warning2;

                    emerg_stop <= 1'b0;
                end
                stop: begin
                    if (((((cur_spd3 == 1'b0) & (cur_spd2 == 1'b0)) & (cur_spd1 == 1'b0)) & (cur_spd0 == 1'b0)))
                        reg_fstate <= stable;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stop;

                    emerg_stop <= 1'b1;
                end
                default: begin
                    emerg_stop <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // speed_control_sm
