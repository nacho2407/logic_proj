// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Mon Dec 23 21:01:46 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module door_open_beep (
    input wire reset,
    input wire clock,
    input wire tick4,
    output reg en,
    output reg [9:0] piano
	 );
	 
    reg [20:0] fstate;
    reg [20:0] reg_fstate;
    localparam n_c12=0,n_n13=1,n_c14=2,n_c15=3,n_n16=4,n_start=5,n_set=6,n_c1=7,n_g2=8,n_e3=9,n_g4=10,n_c5=11,n_c6=12,n_n7=13,n_n8=14,n_n9=15,n_n10=16,n_c11=17,n_ready=18,n_c17=19,n_c18=20;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or tick4)
    begin
        if (reset) begin
            reg_fstate <= n_start;
            en <= 1'b0;
            piano <= 10'b0000000000;
        end
        else begin
            en <= 1'b0;
            piano <= 10'b0000000000;
            case (fstate)
                n_c12: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n13;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c12;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_n13: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n13;

                    en <= 1'b0;
                end
                n_c14: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c15;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c14;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_c15: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n16;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c15;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_n16: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c17;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n16;

                    en <= 1'b0;
                end
                n_start: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_set;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_start;

                    en <= 1'b0;
                end
                n_set: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_set;

                    en <= 1'b0;
                end
                n_c1: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c1;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_g2: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_e3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g2;

                    piano <= 10'b0100000000;

                    en <= 1'b1;
                end
                n_e3: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_e3;

                    piano <= 10'b0001000000;

                    en <= 1'b1;
                end
                n_g4: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g4;

                    piano <= 10'b0100000000;

                    en <= 1'b1;
                end
                n_c5: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c5;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_c6: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c6;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_n7: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n7;

                    en <= 1'b0;
                end
                n_n8: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n8;

                    en <= 1'b0;
                end
                n_n9: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n9;

                    en <= 1'b0;
                end
                n_n10: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c11;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n10;

                    en <= 1'b0;
                end
                n_c11: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c12;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c11;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_ready: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_ready;

                    en <= 1'b0;
                end
                n_c17: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c18;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c17;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_c18: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c18;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                default: begin
                    en <= 1'bx;
                    piano <= 10'bxxxxxxxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // door_open_beep
