// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Sat Dec 21 21:45:54 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module error_beep (
    input wire reset,
    input wire clock,
    input wire tick,
    output reg en,
    output reg [9:0] piano
);

    reg [12:0] fstate;
    reg [12:0] reg_fstate;
    parameter n_start=0,n_set=1,n_m1=2,n_m2=3,n_m3=4,n_m4=5,n_m5=6,n_m6=7,n_m7=8,n_m8=9,n_m9=10,n_m10=11,n_ready=12;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or tick)
    begin
        if (reset) begin
            reg_fstate <= n_start;
            en <= 1'b0;
            piano <= 10'b0000000000;
        end
        else begin
            en <= 1'b0;
            piano <= 10'b0000000000;
            case (fstate)
                n_start: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_set;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_start;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                n_set: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_set;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                n_m1: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m1;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_m2: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m2;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_m3: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m3;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                n_m4: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m4;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                n_m5: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m5;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_m6: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m6;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_m7: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m7;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                n_m8: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m8;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                n_m9: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_m10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m9;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_m10: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_m10;

                    piano <= 10'b1000000000;

                    en <= 1'b1;
                end
                n_ready: begin
                    if ((tick == 1'b1))
                        reg_fstate <= n_ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_ready;

                    piano <= 10'b0000000000;

                    en <= 1'b0;
                end
                default: begin
                    en <= 1'bx;
                    piano <= 10'bxxxxxxxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // error_beep
