// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Mon Dec 23 21:01:46 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module stat_melodyy (
    input wire reset,
    input wire clock,
    input wire tick4,
    output reg en,
    output reg [9:0] piano
	 );
	 
    reg [20:0] fstate;
    reg [20:0] reg_fstate;
    localparam n_start=0, n_set=1, n_c1=2, n_g2=3, n_c3=4, n_d4=5, n_e5=6, n_d6=7, n_c7=8, n_g8=9, n_a9=10, n_f10=11, n_a11=12, n_c12=13, n_f13=14, n_n14=15, n_n15=16, n_n16=17, n_b17=18, n_g18=19, n_b19=20, n_d20=21, n_g21=22, n_f22=23, n_e23=24, n_d24=25, n_e25=26, n_g26=27, n_d27=28, n_g28=29, n_c29=30, n_c30=31, n_ready=32;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or tick4)
    begin
        if (reset) begin
            reg_fstate <= n_start;
            en <= 1'b0;
            piano <= 10'b0000000000;
        end
        else begin
            en <= 1'b0;
            piano <= 10'b0000000000;
            case (fstate)
                n_start: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_set;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_start;

                    en <= 1'b0;
                end
                n_set: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_set;

                    en <= 1'b0;
                end
                n_c1: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c1;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_g2: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g2;

                    piano <= 10'b0000000010;

                    en <= 1'b1;
                end
                n_c3: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_d4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c3;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_d4: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_e5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_d4;

                    piano <= 10'b0000100000;

                    en <= 1'b1;
                end
                n_e5: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_d6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_e5;

                    piano <= 10'b0001000000;

                    en <= 1'b1;
                end
                n_d6: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_d6;

                    piano <= 10'b0000100000;

                    en <= 1'b1;
                end
                n_c7: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c7;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_g8: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_a9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g8;

                    piano <= 10'b0000000010;

                    en <= 1'b1;
                end
                n_a9: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_f10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_a9;

                    piano <= 10'b00000000100;

                    en <= 1'b1;
                end
                n_f10: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_a11;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_f10;

                    piano <= 10'b0000000001;

                    en <= 1'b1;
                end
                n_a11: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c12;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_a11;

                    piano <= 10'b00000000100;

                    en <= 1'b1;
                end
                n_c12: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_f13;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c12;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_f13: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_f13;

                    piano <= 10'b0010000000;

                    en <= 1'b1;
                end
                n_n14: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n15;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n14;

                    en <= 1'b0;
                end
                n_n15: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_n16;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n15;

                    en <= 1'b0;
                end
                n_n16: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_b17;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_n16;

                    en <= 1'b0;
                end
                n_b17: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g18;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_b17;

                    piano <= 10'b0000001000;

                    en <= 1'b1;
                end
                n_g18: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_b19;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g18;

                    piano <= 10'b0000000010;

                    en <= 1'b1;
                end
                n_b19: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_d20;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_b19;

                    piano <= 10'b0000001000;

                    en <= 1'b1;
                end
                n_d20: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g21;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_d20;

                    piano <= 10'b0000100000;

                    en <= 1'b1;
                end
                n_g21: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_f22;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g21;

                    piano <= 10'b0100000000;

                    en <= 1'b1;
                end
                n_f22: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_e23;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_f22;

                    piano <= 10'b0010000000;

                    en <= 1'b1;
                end
                n_e23: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_d24;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_e23;

                    piano <= 10'b0001000000;

                    en <= 1'b1;
                end
					 n_d24: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_e25;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_d24;

                    piano <= 10'b0000100000;

                    en <= 1'b1;
                end
					 n_e25: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g26;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_e25;

                    piano <= 10'b0001000000;

                    en <= 1'b1;
                end
                n_g26: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_d27;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g26;

                    piano <= 10'b0100000000;

                    en <= 1'b1;
                end
					 n_d27: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_g28;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_d27;

                    piano <= 10'b0000100000;

                    en <= 1'b1;
                end
                n_g28: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c29;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_g28;

                    piano <= 10'b0100000000;

                    en <= 1'b1;
                end
                n_c29: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_c30;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c29;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_c30: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_c30;

                    piano <= 10'b0000010000;

                    en <= 1'b1;
                end
                n_ready: begin
                    if ((tick4 == 1'b1))
                        reg_fstate <= n_ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= n_ready;

                    en <= 1'b0;
                end
                default: begin
                    en <= 1'bx;
                    piano <= 10'bxxxxxxxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // stat_melodyy
