// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Fri Dec 13 00:23:51 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module traffic_lt_sm (
    reset,clock,emerg_stop,section_loc3,section_loc0,tik,
    light1,light0,is_stop);

    input reset;
    input clock;
    input emerg_stop;
    input section_loc3;
    input section_loc0;
    input tik;
    tri0 reset;
    tri0 emerg_stop;
    tri0 section_loc3;
    tri0 section_loc0;
    tri0 tik;
    output light1;
    output light0;
    output is_stop;
    reg light1;
    reg light0;
    reg is_stop;
    reg [6:0] fstate;
    reg [6:0] reg_fstate;
    parameter stop=0,wait1=1,wait2=2,ready=3,run=4,stop_ready=5,force_stop=6;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or emerg_stop or section_loc3 or section_loc0 or tik)
    begin
        if (reset) begin
            reg_fstate <= stop;
            light1 <= 1'b0;
            light0 <= 1'b0;
            is_stop <= 1'b0;
        end
        else begin
            light1 <= 1'b0;
            light0 <= 1'b0;
            is_stop <= 1'b0;
            case (fstate)
                stop: begin
                    if (((emerg_stop != 1'b1) & (tik == 1'b1)))
                        reg_fstate <= wait1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stop;

                    is_stop <= 1'b1;

                    light0 <= 1'b1;

                    light1 <= 1'b0;
                end
                wait1: begin
                    if (((emerg_stop != 1'b1) & (tik == 1'b1)))
                        reg_fstate <= wait2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= wait1;

                    is_stop <= 1'b0;

                    light0 <= 1'b1;

                    light1 <= 1'b0;
                end
                wait2: begin
                    if (((emerg_stop != 1'b1) & (tik == 1'b1)))
                        reg_fstate <= ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= wait2;

                    is_stop <= 1'b0;

                    light0 <= 1'b1;

                    light1 <= 1'b0;
                end
                ready: begin
                    if (((emerg_stop != 1'b1) & (tik == 1'b1)))
                        reg_fstate <= run;
                    else if ((emerg_stop == 1'b1))
                        reg_fstate <= force_stop;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= ready;

                    is_stop <= 1'b0;

                    light0 <= 1'b0;

                    light1 <= 1'b1;
                end
                run: begin
                    if (((emerg_stop != 1'b1) & (section_loc3 == 1'b1)))
                        reg_fstate <= stop_ready;
                    else if ((emerg_stop == 1'b1))
                        reg_fstate <= force_stop;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= run;

                    is_stop <= 1'b0;

                    light0 <= 1'b1;

                    light1 <= 1'b1;
                end
                stop_ready: begin
                    if (((emerg_stop != 1'b1) & (section_loc0 == 1'b1)))
                        reg_fstate <= stop;
                    else if ((emerg_stop == 1'b1))
                        reg_fstate <= force_stop;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stop_ready;

                    is_stop <= 1'b0;

                    light0 <= 1'b0;

                    light1 <= 1'b1;
                end
                force_stop: begin
                    if ((emerg_stop != 1'b1))
                        reg_fstate <= ready;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= force_stop;

                    is_stop <= 1'b0;

                    light0 <= 1'b1;

                    light1 <= 1'b0;
                end
                default: begin
                    light1 <= 1'bx;
                    light0 <= 1'bx;
                    is_stop <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // traffic_lt_sm
