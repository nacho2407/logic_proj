// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Sun Dec 22 22:42:07 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module new_location_sm (reset, clock, section_loc, total_loc_wire, states_wire);
	 
	 input wire reset;
    input wire clock;
    input wire [3:0] section_loc;
    output wire [5:0] total_loc_wire;
    output wire [3:0] states_wire;

	 reg [5:0] total_loc;
    reg [3:0] states;
    reg [10:0] fstate;
    reg [10:0] reg_fstate;
    localparam st1=0,tt1=1,st2=2,tt2=3,st3=4,tt3=5,st4=6,tt4=7,st5=8,tt5=9,st6=10;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or section_loc)
    begin
        if (reset) begin
            reg_fstate <= st1;
            total_loc <= 6'b000000;
            states <= 4'b0000;
        end
        else begin
            total_loc <= 6'b000000;
            states <= 4'b0000;
            case (fstate)
                st1: begin
                    if ((section_loc[3:0] == 4'b0010))
                        reg_fstate <= tt1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st1;

                    states <= 4'b0001;

                    total_loc <= 6'b000001;
                end
                tt1: begin
                    if ((section_loc[3:0] == 4'b0001))
                        reg_fstate <= st2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= tt1;

                    states <= 4'b0010;

                    total_loc <= 6'b000001;
                end
                st2: begin
                    if ((section_loc[3:0] == 4'b0010))
                        reg_fstate <= tt2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st2;

                    states <= 4'b0100;

                    total_loc <= 6'b000010;
                end
                tt2: begin
                    if ((section_loc[3:0] == 4'b0001))
                        reg_fstate <= st3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= tt2;

                    states <= 4'b1000;

                    total_loc <= 6'b000010;
                end
                st3: begin
                    if ((section_loc[3:0] == 4'b0010))
                        reg_fstate <= tt3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st3;

                    states <= 4'b0000;

                    total_loc <= 6'b000100;
                end
                tt3: begin
                    if ((section_loc[3:0] == 4'b0001))
                        reg_fstate <= st4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= tt3;

                    states <= 4'b0000;

                    total_loc <= 6'b000100;
                end
                st4: begin
                    if ((section_loc[3:0] == 4'b0010))
                        reg_fstate <= tt4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st4;

                    states <= 4'b0000;

                    total_loc <= 6'b001000;
                end
                tt4: begin
                    if ((section_loc[3:0] == 4'b0001))
                        reg_fstate <= st5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= tt4;

                    states <= 4'b0000;

                    total_loc <= 6'b001000;
                end
                st5: begin
                    if ((section_loc[3:0] == 4'b0010))
                        reg_fstate <= tt5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st5;

                    states <= 4'b0000;

                    total_loc <= 6'b010000;
                end
                tt5: begin
                    if ((section_loc[3:0] == 4'b0001))
                        reg_fstate <= st6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= tt5;

                    states <= 4'b0000;

                    total_loc <= 6'b010000;
                end
                st6: begin
                    if ((section_loc[3:0] == 4'b0010))
                        reg_fstate <= st6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= st6;

                    states <= 4'b0000;

                    total_loc <= 6'b100000;
                end
                default: begin
                    total_loc <= 6'bxxxxxx;
                    states <= 4'bxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // new_location_sm
