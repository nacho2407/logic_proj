// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Sat Dec 14 18:24:50 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module location_sm (
    reset,clock,station1,station0,
    out_tick);

    input reset;
    input clock;
    input station1;
    input station0;
    tri0 reset;
    tri0 station1;
    tri0 station0;
    output out_tick;
    reg out_tick;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter init=0,stable=1,up=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or station1 or station0)
    begin
        if (reset) begin
            reg_fstate <= init;
            out_tick <= 1'b0;
        end
        else begin
            out_tick <= 1'b0;
            case (fstate)
                init: begin
                    if ((station1 == 1'b1))
                        reg_fstate <= stable;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= init;

                    out_tick <= 1'b0;
                end
                stable: begin
                    if ((station0 == 1'b1))
                        reg_fstate <= up;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= stable;

                    out_tick <= 1'b0;
                end
                up: begin
                    if ((station0 == 1'b0))
                        reg_fstate <= stable;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= up;

                    out_tick <= 1'b1;
                end
                default: begin
                    out_tick <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // location_sm
